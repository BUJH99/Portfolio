/********************************************************************************
*
* Module: clock_enable_generator
*
* Description:
*   100MHz의 시스템 클럭(iClk)을 입력받아 6.25MHz 주파수에 해당하는
*   클럭 인에이블(o_wEnClk) 신호를 생성합니다.
*
********************************************************************************/
module clock_enable_generator (
    //==================================================================
    // Port Declarations
    //==================================================================
    input  wire         iClk,       // 시스템 클럭 입력 (100MHz)
    input  wire         iRst_n,       // 시스템 리셋 (active-low)
    output wire         o_wEnClk    // 클럭 인에이블 출력 (6.25MHz 펄스)
);

    //==================================================================
    // Internal Counter Register
    //==================================================================
    // 16분주를 위해 0부터 15까지 카운트하는 4비트 레지스터 (2^4 = 16)
    reg [3:0] count_reg;

    //==================================================================
    // Sequential Logic: Counter
    //==================================================================
    // 시스템 클럭의 상승 엣지마다 카운터를 1씩 증가시킵니다.
    always @(posedge iClk or negedge iRst_n) begin
        if (!iRst_n) begin
            // 시스템 리셋 시, 카운터를 0으로 초기화합니다.
            count_reg <= 4'b0;
        end else begin
            // 카운터가 최대값(15)에 도달하면 0으로 롤오버(Roll-over)합니다.
            if (count_reg == 4'd15) begin
                count_reg <= 4'b0;
            end else begin
                // 그 외의 경우, 카운터를 1 증가시킵니다.
                count_reg <= count_reg + 1'b1;
            end
        end
    end

    //==================================================================
    // Combinational Logic: Output Generation
    //==================================================================
    // 카운터 값이 최대값(15)일 때만 출력 신호를 1로 설정합니다.
    // 이는 정확히 16 클럭마다 한 번씩 발생하는, 1 클럭 폭의 인에이블 펄스를 생성합니다.
    assign o_wEnClk = (count_reg == 4'd15);

endmodule